#############################################################################################
#
#	Copyright 2014-2020 Siemens Product Lifecycle Management Software Inc.
#				All Rights Reserved.
#
#############################################################################################

MACHINE SINUMERIK

EVENT auxfun
{
   UI_LABEL "Auxfun"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM auxfun
   {
      TYPE   i
      DEFVAL "0"
      UI_LABEL "Auxfun Value"
   }
   PARAM auxfun_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT coolant_off
{
   UI_LABEL "Coolant Off"
   CATEGORY MILL DRILL LATHE

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM coolant_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT set_pocket4_parameters
{
   UI_LABEL "Set POCKET4 Parameters"
   CATEGORY MILL DRILL

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM pocket4_maximum_infeed_width
   {
      TYPE   d
      DEFVAL "0.0000"
      UI_LABEL "Maximum Infeed Width"
   }
   PARAM pocket4_helical_path_radius
   {
      TYPE   d
      DEFVAL "2.0000"
      UI_LABEL "Helical Path Radius"
   }
}

EVENT dwell
{
   POST_EVENT "delay"
   UI_LABEL "Dwell"

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM delay_mode
   {
      TYPE o
      DEFVAL "Seconds"
      OPTIONS "Seconds","Revolutions"
      UI_LABEL "Dwell Type"
   }
   PARAM delay_value
   {
      TYPE   d
      DEFVAL "10.0000"
      UI_LABEL "Dwell Value"
   }
   PARAM delay_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT insert
{
   UI_LABEL "Insert"

   PARAM Instruction
   {
      TYPE    s
   }
}

EVENT length_compensation
{
   UI_LABEL "Tool Length Compensation"
   CATEGORY MILL DRILL LATHE

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM Overide_operation_param
   {
      TYPE   b
      DEFVAL "TRUE"
      UI_LABEL "Override Operation Parameter"
   }
   PARAM length_comp_register
   {
      TYPE   i
      DEFVAL "2"
      UI_LABEL "Adjust Register"
   }
   PARAM length_comp_register_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT opskip_on
{
   UI_LABEL "Optional Skip On"

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM opskip_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT opskip_off
{
   UI_LABEL "Optional Skip Off"

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM opskip_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT opstop
{
   UI_LABEL "Optional Stop"

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM opstop_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT prefer_solution
{
	UI_LABEL "Preferred Solution"
	PARAM command_status
	{
		TYPE o
		DEFVAL "Active"
		OPTIONS "Active","Inactive","User Defined"
		UI_LABEL "Status"
	}
	PARAM prefer_axis
	{
		TYPE o
		DEFVAL "OFF"
		OPTIONS "OFF", "A", "B", "C"
		UI_LABEL "Preferred Axis"
	}
	PARAM prefer_output_min
	{
		TYPE d
		DEFVAL "0.000000"
		TOGGLE Off
		UI_LABEL "Preferred Range Minimum"
	}
	PARAM prefer_output_max
	{
		TYPE d
		DEFVAL "0.000000"
		TOGGLE Off
		UI_LABEL "Preferred Range Maximum"
	}
}


EVENT prefun
{
   UI_LABEL "Prefun"

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM prefun
   {
      TYPE   i
      DEFVAL "0"
      UI_LABEL "Prefun Value"
   }
   PARAM prefun_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT rotate
{
   UI_LABEL "Rotate"
   CATEGORY MILL DRILL LATHE

   PARAM command_status
   {
      TYPE o
      DEFVAL   "Active"
      OPTIONS  "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM rotate_axis_type
   {
      TYPE o
      DEFVAL   "Table"
      OPTIONS  "Table","Head","Aaxis","Baxis","Caxis","Fourth_Axis","Fifth_Axis"
      UI_LABEL "Rotation Axis"
   }
   PARAM rotation_mode
   {
      TYPE o
      DEFVAL   "None"
      OPTIONS  "None","Angle","Absolute","Incremental"
      UI_LABEL "Type"
   }
   PARAM rotation_direction
   {
      TYPE   o
      DEFVAL   "CLW"
      OPTIONS  "CLW","CCLW","NONE"
      UI_LABEL "Direction"
   }
   PARAM rotation_angle
   {
      TYPE   d
      DEFVAL   "0.0000"
      TOGGLE   On
      UI_LABEL "Angle"
   }
   PARAM rotation_reference_mode
   {
      TYPE   b
      DEFVAL "FALSE"
      UI_LABEL "Reference Only - No Output"
   }
   PARAM rotation_text
   {
      TYPE   s
      TOGGLE   Off
      UI_LABEL "Text"
   }
}

EVENT sequence_number
{
   UI_LABEL "Sequence Number"

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM sequence_mode
   {
      TYPE o
      DEFVAL "N"
      OPTIONS "N","Off","On","Auto"
      UI_LABEL "Number Type"
   }
   PARAM sequence_number
   {
      TYPE   i
      DEFVAL "0"
      UI_LABEL "Number"
   }
   PARAM sequence_increment
   {
      TYPE   i
      DEFVAL "0"
      UI_LABEL "Increment"
   }
   PARAM sequence_frequency
   {
      TYPE   i
      DEFVAL "0"
      UI_LABEL "Frequency"
   }
   PARAM sequence_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT stop
{
   UI_LABEL "Stop"

   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM stop_text
   {
      TYPE   s
      TOGGLE Off
      UI_LABEL "Text"
   }
}

EVENT text
{
   UI_LABEL "User Defined"

   PARAM user_defined_text
   {
      TYPE   s
      TOGGLE On
      UI_LABEL "User Defined Command"
   }
}

EVENT structure_representation_mode
{
   UI_LABEL "Operation representation in collpased mode"
   PARAM output_status
   {
      TYPE o
      DEFVAL "On"
      OPTIONS "On","Off"
      UI_LABEL "Output"
   }
   PARAM display_name
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Display name"
   }
   PARAM readonly_status
   {
      TYPE o
      DEFVAL "Editable"
      OPTIONS "Editable","Readonly"
      UI_LABEL "Status"
   }
   PARAM type_status
   {
      TYPE o
      DEFVAL "Operation"
      OPTIONS "Header","Operation"
      UI_LABEL "Status"
   }
}

EVENT LIB_manual_CYCLE800_setting
{
   UI_LABEL "Manual CYCLE800 setting"
   PARAM lib_cycle800_dir
   {
      TYPE o
      DEFVAL "Auto"
      OPTIONS "Auto","+1","-1"
      UI_LABEL "Direction"
   }
}

EVENT program_control
{
	UI_LABEL "Program Control"
	CATEGORY MILL DRILL
	PARAM ctrl_program_control
	{
		TYPE b
		DEFVAL "FALSE"
		UI_LABEL "Call External Subroutine for Each Operation"
	}
}
